module lab9_3(HEX0, HEX1, HEX2, HEX3, LEDR, SW, KEY);
	input [9:0] SW;
	input [0:0] KEY;
	output [6:0] HEX0, HEX1, HEX2, HEX3;
	output [0:0] LEDR;

	wire [3:0] out;
	

	ram(SW[8:4], SW[3:0], KEY[0], SW[9], out);
	converter(HEX0, out);
	converter(HEX1, SW[3:0]);
	converter(HEX2, SW[7:4]);
	converter(HEX3, SW[8]);
	
	assign LEDR[0] = SW[9];
endmodule

module ram(address, data, clock, wren, q);
	input [4:0] address;
	input [3:0] data;
	input clock, wren;
	output reg [3:0] q;
	reg [3:0] array[31:0];	
	always @ (posedge clock) begin
		if(wren)
			array[address] <= data;
	
		q <= array[address];
	end
endmodule

module converter(seg, num);
	 input [3:0] num;
	 output reg [6:0] seg;
    always @(num) begin
        case (num)
			4'b0000: seg <= 7'b1000000; // 0
			4'b0001: seg <= 7'b1111001; // 1
			4'b0010: seg <= 7'b0100100; // 2
			4'b0011: seg <= 7'b0110000; // 3
			4'b0100: seg <= 7'b0011001; // 4
			4'b0101: seg <= 7'b0010010; // 5
			4'b0110: seg <= 7'b0000010; // 6
			4'b0111: seg <= 7'b1111000; // 7
			4'b1000: seg <= 7'b0000000; // 8
			4'b1001: seg <= 7'b0011000; // 9
			4'b1010: seg <= 7'b0001000; // A
			4'b1011: seg <= 7'b0000000; // B
			4'b1100: seg <= 7'b1000110; // C
			4'b1101: seg <= 7'b1000000; // D
			4'b1110: seg <= 7'b0000110; // E
			4'b1111: seg <= 7'b0001110; // F
			default: seg <= 7'b0000000; //  
       endcase
    end
endmodule